`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module BranchAdd(
    input [31:0] ShiftLeft2,
    input [31:0] PCAdd,
    output [31:0] BranchAddOut

    );
    assign BranchAddOut = ShiftLeft2+PCAdd;
endmodule
